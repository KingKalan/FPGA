// Placeholder top-level module
module numen_top(); endmodule
